-------------------------------------------------------------------------------
--                                                                      
--                        4x7-segments counter project
--  
-------------------------------------------------------------------------------
--                                                                      
--
-- FILENAME:                io_ctrl_rtl.vhd
-- 
-- ENGINEER:                Moritz Emersberger
--  
-- DATE (current Version):  31. March 2023
--  
-- VERSION:                 1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION: The IO Control unit is part of the counter project.
--              It manages the interface to the 7-segment displays,
--              the LEDs, the push buttons and the switches of the
--              Digilent Basys3 FPGA board   
--
-------------------------------------------------------------------------------
--                                                                      
-- CHANGES:     V1.0: 31.03.2023: initial Version     
--
-------------------------------------------------------------------------------

configuration io_ctrl_rtl_cfg of io_ctrl is
  for rtl        
  end for;
end io_ctrl_rtl_cfg;
